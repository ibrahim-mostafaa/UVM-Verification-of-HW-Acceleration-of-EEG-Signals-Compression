`include "uvm_pkg.sv"

package pack1;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "Seq_Item.sv"
	`include "Sequence.sv"
	`include "Sequencer.sv"
	`include "Driver.sv"
	`include "Monitor.sv"
	`include "Scoreboard.sv"
	`include "Subscriber.sv"
	`include "Agent.sv"
	`include "Env.sv"
	`include "Test.sv"
endpackage : pack1


